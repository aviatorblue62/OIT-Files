// <Houston & Fawver, EE 133 Lab 9 Traffic Light, 05-27-2014>

module traffic_light(
		input wire clk,reset,sensor,
		output reg hwy